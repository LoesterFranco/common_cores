`define ACCESS_PACKED(idx, len) (len)*(idx) +: len